    .tl_CORE_NAME_scratchpad_instr_o(CORE_NAME_scratchpad_instr_req),
    .tl_CORE_NAME_scratchpad_instr_i(CORE_NAME_scratchpad_instr_rsp),
    .tl_CORE_NAME_scratchpad_data_o (CORE_NAME_scratchpad_data_req),
    .tl_CORE_NAME_scratchpad_data_i (CORE_NAME_scratchpad_data_rsp),
