// Copyright (c) 2025 Ben Krusekamp
// Licensed under the Solderpad Hardware License v2.1. See LICENSE file in the project root for details.
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1

tlul_pkg::tl_h2d_t CORE_NAME_scratchpad_instr_req;
tlul_pkg::tl_d2h_t CORE_NAME_scratchpad_instr_rsp;
tlul_pkg::tl_h2d_t CORE_NAME_scratchpad_data_req;
tlul_pkg::tl_d2h_t CORE_NAME_scratchpad_data_rsp;

tlul_pkg::tl_h2d_t CORE_NAME_core_instr_req;
tlul_pkg::tl_d2h_t CORE_NAME_core_instr_rsp;
tlul_pkg::tl_h2d_t CORE_NAME_core_data_req;
tlul_pkg::tl_d2h_t CORE_NAME_core_data_rsp;
