// Copyright (c) 2025 Ben Krusekamp
// Licensed under the Solderpad Hardware License v2.1. See LICENSE file in the project root for details.
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1

    .tl_CORE_NAME_scratchpad_instr_o(CORE_NAME_scratchpad_instr_req),
    .tl_CORE_NAME_scratchpad_instr_i(CORE_NAME_scratchpad_instr_rsp),
    .tl_CORE_NAME_scratchpad_data_o (CORE_NAME_scratchpad_data_req),
    .tl_CORE_NAME_scratchpad_data_i (CORE_NAME_scratchpad_data_rsp),
