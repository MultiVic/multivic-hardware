tlul_pkg::tl_h2d_t CORE_NAME_scratchpad_instr_req;
tlul_pkg::tl_d2h_t CORE_NAME_scratchpad_instr_rsp;
tlul_pkg::tl_h2d_t CORE_NAME_scratchpad_data_req;
tlul_pkg::tl_d2h_t CORE_NAME_scratchpad_data_rsp;

tlul_pkg::tl_h2d_t CORE_NAME_core_instr_req;
tlul_pkg::tl_d2h_t CORE_NAME_core_instr_rsp;
tlul_pkg::tl_h2d_t CORE_NAME_core_data_req;
tlul_pkg::tl_d2h_t CORE_NAME_core_data_rsp;
